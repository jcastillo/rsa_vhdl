--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   17:40:28 12/13/2009
-- Design Name:   
-- Module Name:   C:/ise_wp/ciosspartan/test_rsa_1024.vhd
-- Project Name:  ciosspartan
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: rsa_top
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;
 
ENTITY test_rsa_4096 IS
END test_rsa_4096;
 
ARCHITECTURE behavior OF test_rsa_4096 IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT rsa_top
    PORT(
         clk : IN  std_logic;
         reset : IN  std_logic;
         valid_in : IN  std_logic;
         x : IN  std_logic_vector(15 downto 0);
         y : IN  std_logic_vector(15 downto 0);
         m : IN  std_logic_vector(15 downto 0);
         r_c : IN  std_logic_vector(15 downto 0);
         n_c : IN  std_logic_vector(15 downto 0);
         s : OUT  std_logic_vector(15 downto 0);
         valid_out : OUT  std_logic;
         word_number : IN  std_logic_vector(15 downto 0);
			bit_size : in std_logic_vector(15 downto 0) 
        );
    END COMPONENT;
    
    

   --Inputs
   signal clk : std_logic := '0';
   signal reset : std_logic := '0';
   signal valid_in : std_logic := '0';
   signal x : std_logic_vector(15 downto 0) := (others => '0');
   signal y : std_logic_vector(15 downto 0) := (others => '0');
   signal m : std_logic_vector(15 downto 0) := (others => '0');
   signal r_c : std_logic_vector(15 downto 0) := (others => '0');
   signal n_c : std_logic_vector(15 downto 0) := (others => '0');
   signal word_number : std_logic_vector(15 downto 0) := x"0100";
   signal bit_size : std_logic_vector(15 downto 0) := x"1000";
 	--Outputs
   signal s : std_logic_vector(15 downto 0);
   signal valid_out : std_logic;

   -- Clock period definitions
   constant clk_period : time := 1ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: rsa_top PORT MAP (
          clk => clk,
          reset => reset,
          valid_in => valid_in,
          x => x,
          y => y,
          m => m,
          r_c => r_c,
          n_c => n_c,
          s => s,
          valid_out => valid_out,
          word_number => word_number,
			 bit_size => bit_size
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
	   valid_in<='0';
      -- hold reset state for 100ms.
		reset <= '1';
      wait for 10ns;	
      reset <= '0';
      wait for clk_period*10;

      -- insert stimulus here 

--n_c and valid signal and the r_c constant are also required
		n_c <= x"e5a7";
		valid_in <= '1';
		x <= x"f3ad";
		y <= x"f9e3";
		m <= x"8de9";
		r_c <= x"6f2e";
		wait for clk_period;
		x <= x"8e40";
		y <= x"b134";
		m <= x"d218";
		r_c <= x"6999";
		wait for clk_period;
		x <= x"6af9";
		y <= x"fa23";
		m <= x"3113";
		r_c <= x"77ad";
		wait for clk_period;
		x <= x"4e63";
		y <= x"2b9e";
		m <= x"df1f";
		r_c <= x"d4fd";
		wait for clk_period;
		x <= x"9600";
		y <= x"071b";
		m <= x"6757";
		r_c <= x"44a8";
		wait for clk_period;
		x <= x"68f4";
		y <= x"cfe8";
		m <= x"bc83";
		r_c <= x"95dd";
		wait for clk_period;
		x <= x"5a12";
		y <= x"e5dc";
		m <= x"4bd4";
		r_c <= x"d1c0";
		wait for clk_period;
		x <= x"d62e";
		y <= x"8165";
		m <= x"0eda";
		r_c <= x"06ac";
		wait for clk_period;
		x <= x"8fc1";
		y <= x"5ddc";
		m <= x"18cc";
		r_c <= x"0378";
		wait for clk_period;
		x <= x"d2cd";
		y <= x"12c2";
		m <= x"4b5e";
		r_c <= x"7c54";
		wait for clk_period;
		x <= x"c6e4";
		y <= x"2247";
		m <= x"8233";
		r_c <= x"bce5";
		wait for clk_period;
		x <= x"4a36";
		y <= x"361f";
		m <= x"3ff4";
		r_c <= x"379f";
		wait for clk_period;
		x <= x"cedf";
		y <= x"13c6";
		m <= x"fdf8";
		r_c <= x"cf64";
		wait for clk_period;
		x <= x"19ea";
		y <= x"a4a6";
		m <= x"add6";
		r_c <= x"960f";
		wait for clk_period;
		x <= x"ad18";
		y <= x"3ce3";
		m <= x"8a5c";
		r_c <= x"a637";
		wait for clk_period;
		x <= x"4402";
		y <= x"b6cf";
		m <= x"7112";
		r_c <= x"f8aa";
		wait for clk_period;
		x <= x"fdb2";
		y <= x"e4b5";
		m <= x"f09b";
		r_c <= x"15af";
		wait for clk_period;
		x <= x"45fa";
		y <= x"6e5c";
		m <= x"2b15";
		r_c <= x"60b0";
		wait for clk_period;
		x <= x"6941";
		y <= x"0e2f";
		m <= x"5ed4";
		r_c <= x"72c0";
		wait for clk_period;
		x <= x"61cf";
		y <= x"7bbd";
		m <= x"1e22";
		r_c <= x"ffad";
		wait for clk_period;
		x <= x"6c80";
		y <= x"4f5a";
		m <= x"f036";
		r_c <= x"c57d";
		wait for clk_period;
		x <= x"2e3c";
		y <= x"b06b";
		m <= x"9968";
		r_c <= x"8944";
		wait for clk_period;
		x <= x"b5c5";
		y <= x"4871";
		m <= x"07fd";
		r_c <= x"2775";
		wait for clk_period;
		x <= x"f44b";
		y <= x"056d";
		m <= x"8b1a";
		r_c <= x"d40e";
		wait for clk_period;
		x <= x"f9c6";
		y <= x"50aa";
		m <= x"0e08";
		r_c <= x"23af";
		wait for clk_period;
		x <= x"e9a2";
		y <= x"4881";
		m <= x"3eb2";
		r_c <= x"2d22";
		wait for clk_period;
		x <= x"2148";
		y <= x"b560";
		m <= x"0dbd";
		r_c <= x"69b8";
		wait for clk_period;
		x <= x"b16b";
		y <= x"4a88";
		m <= x"c5d6";
		r_c <= x"ce78";
		wait for clk_period;
		x <= x"4038";
		y <= x"b2e4";
		m <= x"87a5";
		r_c <= x"a4c1";
		wait for clk_period;
		x <= x"4496";
		y <= x"7d58";
		m <= x"6de3";
		r_c <= x"488c";
		wait for clk_period;
		x <= x"99f0";
		y <= x"8d9b";
		m <= x"a222";
		r_c <= x"8f06";
		wait for clk_period;
		x <= x"7560";
		y <= x"6815";
		m <= x"4998";
		r_c <= x"3a95";
		wait for clk_period;
		x <= x"9fe3";
		y <= x"d930";
		m <= x"726c";
		r_c <= x"54a1";
		wait for clk_period;
		x <= x"5579";
		y <= x"39c2";
		m <= x"918c";
		r_c <= x"4e47";
		wait for clk_period;
		x <= x"74b5";
		y <= x"affb";
		m <= x"fc29";
		r_c <= x"963f";
		wait for clk_period;
		x <= x"71e4";
		y <= x"a485";
		m <= x"627c";
		r_c <= x"1b4c";
		wait for clk_period;
		x <= x"45e6";
		y <= x"7d24";
		m <= x"6ffc";
		r_c <= x"1bee";
		wait for clk_period;
		x <= x"f595";
		y <= x"2205";
		m <= x"9778";
		r_c <= x"fb33";
		wait for clk_period;
		x <= x"91e3";
		y <= x"f457";
		m <= x"307a";
		r_c <= x"e5fc";
		wait for clk_period;
		x <= x"4ef1";
		y <= x"1e9d";
		m <= x"86e4";
		r_c <= x"beff";
		wait for clk_period;
		x <= x"d694";
		y <= x"692c";
		m <= x"3e46";
		r_c <= x"f818";
		wait for clk_period;
		x <= x"475c";
		y <= x"ee38";
		m <= x"1866";
		r_c <= x"fae5";
		wait for clk_period;
		x <= x"9b2b";
		y <= x"8b0d";
		m <= x"f740";
		r_c <= x"9921";
		wait for clk_period;
		x <= x"e3fc";
		y <= x"a94c";
		m <= x"143d";
		r_c <= x"8503";
		wait for clk_period;
		x <= x"2009";
		y <= x"9da9";
		m <= x"a1d5";
		r_c <= x"b9ba";
		wait for clk_period;
		x <= x"2aa1";
		y <= x"4350";
		m <= x"ac64";
		r_c <= x"92ad";
		wait for clk_period;
		x <= x"9f13";
		y <= x"8d5c";
		m <= x"c532";
		r_c <= x"fa04";
		wait for clk_period;
		x <= x"6672";
		y <= x"160d";
		m <= x"cc81";
		r_c <= x"363e";
		wait for clk_period;
		x <= x"f315";
		y <= x"19f9";
		m <= x"fda1";
		r_c <= x"4fd5";
		wait for clk_period;
		x <= x"adf5";
		y <= x"0fc9";
		m <= x"0b5e";
		r_c <= x"5ca7";
		wait for clk_period;
		x <= x"5c95";
		y <= x"e8ac";
		m <= x"9f10";
		r_c <= x"95a2";
		wait for clk_period;
		x <= x"228f";
		y <= x"7096";
		m <= x"24b6";
		r_c <= x"6408";
		wait for clk_period;
		x <= x"f2d3";
		y <= x"6f97";
		m <= x"171d";
		r_c <= x"00e6";
		wait for clk_period;
		x <= x"2306";
		y <= x"3906";
		m <= x"8a04";
		r_c <= x"7d8f";
		wait for clk_period;
		x <= x"e5e0";
		y <= x"821b";
		m <= x"a882";
		r_c <= x"df3d";
		wait for clk_period;
		x <= x"93b7";
		y <= x"69fd";
		m <= x"481a";
		r_c <= x"5b5b";
		wait for clk_period;
		x <= x"1f17";
		y <= x"389c";
		m <= x"8df8";
		r_c <= x"3623";
		wait for clk_period;
		x <= x"48fd";
		y <= x"459d";
		m <= x"d75e";
		r_c <= x"43ea";
		wait for clk_period;
		x <= x"257f";
		y <= x"e6b0";
		m <= x"f557";
		r_c <= x"ff2e";
		wait for clk_period;
		x <= x"b9f2";
		y <= x"4d40";
		m <= x"e983";
		r_c <= x"6f0c";
		wait for clk_period;
		x <= x"4e80";
		y <= x"2568";
		m <= x"e60b";
		r_c <= x"2cd6";
		wait for clk_period;
		x <= x"698f";
		y <= x"5539";
		m <= x"f50f";
		r_c <= x"06d3";
		wait for clk_period;
		x <= x"fccb";
		y <= x"e6cc";
		m <= x"719c";
		r_c <= x"b995";
		wait for clk_period;
		x <= x"3adc";
		y <= x"bbc9";
		m <= x"b749";
		r_c <= x"8604";
		wait for clk_period;
		x <= x"e40f";
		y <= x"2136";
		m <= x"50cf";
		r_c <= x"3b02";
		wait for clk_period;
		x <= x"af98";
		y <= x"b1e0";
		m <= x"fb9c";
		r_c <= x"7bf6";
		wait for clk_period;
		x <= x"e636";
		y <= x"cab6";
		m <= x"c8db";
		r_c <= x"8be7";
		wait for clk_period;
		x <= x"6004";
		y <= x"fd63";
		m <= x"d65b";
		r_c <= x"5c90";
		wait for clk_period;
		x <= x"8f49";
		y <= x"8d5c";
		m <= x"a390";
		r_c <= x"8c07";
		wait for clk_period;
		x <= x"a126";
		y <= x"4baf";
		m <= x"345d";
		r_c <= x"309f";
		wait for clk_period;
		x <= x"62e5";
		y <= x"2e2d";
		m <= x"7f9b";
		r_c <= x"204c";
		wait for clk_period;
		x <= x"fc1d";
		y <= x"b6d7";
		m <= x"af98";
		r_c <= x"32e2";
		wait for clk_period;
		x <= x"2cd8";
		y <= x"6c1d";
		m <= x"c18c";
		r_c <= x"fbcf";
		wait for clk_period;
		x <= x"6e4d";
		y <= x"c04f";
		m <= x"a645";
		r_c <= x"c45d";
		wait for clk_period;
		x <= x"a36c";
		y <= x"f1df";
		m <= x"e409";
		r_c <= x"0c8c";
		wait for clk_period;
		x <= x"edf4";
		y <= x"9216";
		m <= x"ace6";
		r_c <= x"74f6";
		wait for clk_period;
		x <= x"9eac";
		y <= x"cdbe";
		m <= x"cfce";
		r_c <= x"db6b";
		wait for clk_period;
		x <= x"d181";
		y <= x"2d49";
		m <= x"dc88";
		r_c <= x"ae65";
		wait for clk_period;
		x <= x"402a";
		y <= x"7dc6";
		m <= x"9318";
		r_c <= x"abc0";
		wait for clk_period;
		x <= x"db24";
		y <= x"c31f";
		m <= x"e05b";
		r_c <= x"d176";
		wait for clk_period;
		x <= x"5faf";
		y <= x"0065";
		m <= x"3278";
		r_c <= x"5916";
		wait for clk_period;
		x <= x"9414";
		y <= x"d5a1";
		m <= x"514d";
		r_c <= x"3dea";
		wait for clk_period;
		x <= x"1cf6";
		y <= x"5c21";
		m <= x"074a";
		r_c <= x"7e1c";
		wait for clk_period;
		x <= x"c806";
		y <= x"a8ff";
		m <= x"1eee";
		r_c <= x"9ec4";
		wait for clk_period;
		x <= x"e3c6";
		y <= x"f7c8";
		m <= x"c5fd";
		r_c <= x"27e5";
		wait for clk_period;
		x <= x"5c52";
		y <= x"0179";
		m <= x"d901";
		r_c <= x"59ba";
		wait for clk_period;
		x <= x"44bb";
		y <= x"2e2d";
		m <= x"c5f1";
		r_c <= x"fdf9";
		wait for clk_period;
		x <= x"9c6f";
		y <= x"8970";
		m <= x"7231";
		r_c <= x"adf5";
		wait for clk_period;
		x <= x"9a2f";
		y <= x"eb49";
		m <= x"938d";
		r_c <= x"cdcb";
		wait for clk_period;
		x <= x"148e";
		y <= x"b741";
		m <= x"348c";
		r_c <= x"bd49";
		wait for clk_period;
		x <= x"16b2";
		y <= x"825b";
		m <= x"5bad";
		r_c <= x"91b8";
		wait for clk_period;
		x <= x"038b";
		y <= x"f0f8";
		m <= x"15ac";
		r_c <= x"fb48";
		wait for clk_period;
		x <= x"4964";
		y <= x"9ece";
		m <= x"0ff4";
		r_c <= x"15c9";
		wait for clk_period;
		x <= x"9f04";
		y <= x"8677";
		m <= x"08d4";
		r_c <= x"b188";
		wait for clk_period;
		x <= x"5609";
		y <= x"4a98";
		m <= x"9b9a";
		r_c <= x"18dd";
		wait for clk_period;
		x <= x"fe37";
		y <= x"baf9";
		m <= x"14a9";
		r_c <= x"e603";
		wait for clk_period;
		x <= x"5799";
		y <= x"24f9";
		m <= x"e1f7";
		r_c <= x"f4f6";
		wait for clk_period;
		x <= x"4b55";
		y <= x"200c";
		m <= x"8d44";
		r_c <= x"b76b";
		wait for clk_period;
		x <= x"1e47";
		y <= x"8e33";
		m <= x"c1ab";
		r_c <= x"0109";
		wait for clk_period;
		x <= x"5e67";
		y <= x"5738";
		m <= x"06bb";
		r_c <= x"82f7";
		wait for clk_period;
		x <= x"5954";
		y <= x"49a0";
		m <= x"3207";
		r_c <= x"fe69";
		wait for clk_period;
		x <= x"1e3f";
		y <= x"8a88";
		m <= x"6f83";
		r_c <= x"0820";
		wait for clk_period;
		x <= x"ef19";
		y <= x"afaf";
		m <= x"a32b";
		r_c <= x"0d81";
		wait for clk_period;
		x <= x"6944";
		y <= x"90e6";
		m <= x"e2a5";
		r_c <= x"444d";
		wait for clk_period;
		x <= x"75cd";
		y <= x"8521";
		m <= x"c8cc";
		r_c <= x"b4d0";
		wait for clk_period;
		x <= x"b2b4";
		y <= x"bd9a";
		m <= x"3254";
		r_c <= x"cece";
		wait for clk_period;
		x <= x"3fc9";
		y <= x"10dc";
		m <= x"0502";
		r_c <= x"51de";
		wait for clk_period;
		x <= x"009e";
		y <= x"5c27";
		m <= x"a76e";
		r_c <= x"b84b";
		wait for clk_period;
		x <= x"87b2";
		y <= x"2109";
		m <= x"b70b";
		r_c <= x"f69f";
		wait for clk_period;
		x <= x"76b9";
		y <= x"7ef4";
		m <= x"e075";
		r_c <= x"a4b8";
		wait for clk_period;
		x <= x"a58a";
		y <= x"d451";
		m <= x"e41d";
		r_c <= x"42c9";
		wait for clk_period;
		x <= x"6a76";
		y <= x"bf83";
		m <= x"5650";
		r_c <= x"2589";
		wait for clk_period;
		x <= x"6a87";
		y <= x"e34c";
		m <= x"1a1e";
		r_c <= x"a367";
		wait for clk_period;
		x <= x"27a8";
		y <= x"a572";
		m <= x"b41b";
		r_c <= x"2a94";
		wait for clk_period;
		x <= x"b198";
		y <= x"9a64";
		m <= x"c014";
		r_c <= x"1c8c";
		wait for clk_period;
		x <= x"1923";
		y <= x"3b82";
		m <= x"6693";
		r_c <= x"1e1f";
		wait for clk_period;
		x <= x"74b0";
		y <= x"70b4";
		m <= x"6c37";
		r_c <= x"0e84";
		wait for clk_period;
		x <= x"c283";
		y <= x"4ca1";
		m <= x"3289";
		r_c <= x"91e1";
		wait for clk_period;
		x <= x"2634";
		y <= x"f221";
		m <= x"85fa";
		r_c <= x"514a";
		wait for clk_period;
		x <= x"7347";
		y <= x"00bf";
		m <= x"9055";
		r_c <= x"bdbc";
		wait for clk_period;
		x <= x"6f26";
		y <= x"f955";
		m <= x"2bc2";
		r_c <= x"b92c";
		wait for clk_period;
		x <= x"6423";
		y <= x"33e4";
		m <= x"feb0";
		r_c <= x"4c60";
		wait for clk_period;
		x <= x"8723";
		y <= x"3393";
		m <= x"3410";
		r_c <= x"81eb";
		wait for clk_period;
		x <= x"7346";
		y <= x"b1e1";
		m <= x"52b0";
		r_c <= x"002d";
		wait for clk_period;
		x <= x"fbc2";
		y <= x"1104";
		m <= x"922b";
		r_c <= x"2801";
		wait for clk_period;
		x <= x"346a";
		y <= x"9a47";
		m <= x"eb77";
		r_c <= x"796d";
		wait for clk_period;
		x <= x"6827";
		y <= x"5712";
		m <= x"7523";
		r_c <= x"38c5";
		wait for clk_period;
		x <= x"8374";
		y <= x"353e";
		m <= x"3843";
		r_c <= x"39e5";
		wait for clk_period;
		x <= x"b9f2";
		y <= x"3458";
		m <= x"ce86";
		r_c <= x"949d";
		wait for clk_period;
		x <= x"4e80";
		y <= x"15b7";
		m <= x"a092";
		r_c <= x"faef";
		wait for clk_period;
		x <= x"698f";
		y <= x"79d3";
		m <= x"b6bc";
		r_c <= x"49bf";
		wait for clk_period;
		x <= x"fccb";
		y <= x"36fa";
		m <= x"d277";
		r_c <= x"7cc1";
		wait for clk_period;
		x <= x"3adc";
		y <= x"b005";
		m <= x"8807";
		r_c <= x"298f";
		wait for clk_period;
		x <= x"e40f";
		y <= x"6417";
		m <= x"9623";
		r_c <= x"a58e";
		wait for clk_period;
		x <= x"af98";
		y <= x"4b5e";
		m <= x"710d";
		r_c <= x"db3c";
		wait for clk_period;
		x <= x"e636";
		y <= x"4312";
		m <= x"e49b";
		r_c <= x"8961";
		wait for clk_period;
		x <= x"6004";
		y <= x"7ee9";
		m <= x"3e5d";
		r_c <= x"9aae";
		wait for clk_period;
		x <= x"8f49";
		y <= x"85bd";
		m <= x"489c";
		r_c <= x"ad8d";
		wait for clk_period;
		x <= x"a126";
		y <= x"fd6b";
		m <= x"fc21";
		r_c <= x"0a91";
		wait for clk_period;
		x <= x"62e5";
		y <= x"0dd3";
		m <= x"14bd";
		r_c <= x"729e";
		wait for clk_period;
		x <= x"fc1d";
		y <= x"e766";
		m <= x"5b19";
		r_c <= x"c082";
		wait for clk_period;
		x <= x"2cd8";
		y <= x"e716";
		m <= x"daa2";
		r_c <= x"2329";
		wait for clk_period;
		x <= x"6e4d";
		y <= x"f905";
		m <= x"f588";
		r_c <= x"4f43";
		wait for clk_period;
		x <= x"a36c";
		y <= x"454f";
		m <= x"67f7";
		r_c <= x"1b0b";
		wait for clk_period;
		x <= x"edf4";
		y <= x"1e4a";
		m <= x"ad6f";
		r_c <= x"b1f9";
		wait for clk_period;
		x <= x"9eac";
		y <= x"bf1d";
		m <= x"1eab";
		r_c <= x"d230";
		wait for clk_period;
		x <= x"d181";
		y <= x"cd80";
		m <= x"3441";
		r_c <= x"10fd";
		wait for clk_period;
		x <= x"402a";
		y <= x"def8";
		m <= x"4e75";
		r_c <= x"da66";
		wait for clk_period;
		x <= x"db24";
		y <= x"d36e";
		m <= x"3d26";
		r_c <= x"98bd";
		wait for clk_period;
		x <= x"5faf";
		y <= x"b582";
		m <= x"9044";
		r_c <= x"8007";
		wait for clk_period;
		x <= x"9414";
		y <= x"f46f";
		m <= x"6ea7";
		r_c <= x"76a6";
		wait for clk_period;
		x <= x"1cf6";
		y <= x"2188";
		m <= x"324d";
		r_c <= x"4b44";
		wait for clk_period;
		x <= x"c806";
		y <= x"36de";
		m <= x"524d";
		r_c <= x"7132";
		wait for clk_period;
		x <= x"e3c6";
		y <= x"9c7c";
		m <= x"6aba";
		r_c <= x"e9d1";
		wait for clk_period;
		x <= x"5c52";
		y <= x"b727";
		m <= x"92bb";
		r_c <= x"24ae";
		wait for clk_period;
		x <= x"44bb";
		y <= x"6acb";
		m <= x"2031";
		r_c <= x"6da3";
		wait for clk_period;
		x <= x"9c6f";
		y <= x"87d9";
		m <= x"cbc6";
		r_c <= x"9d56";
		wait for clk_period;
		x <= x"9a2f";
		y <= x"5cc6";
		m <= x"8b29";
		r_c <= x"f989";
		wait for clk_period;
		x <= x"148e";
		y <= x"e3e4";
		m <= x"55d6";
		r_c <= x"acf9";
		wait for clk_period;
		x <= x"16b2";
		y <= x"496a";
		m <= x"ee20";
		r_c <= x"3203";
		wait for clk_period;
		x <= x"038b";
		y <= x"d3a9";
		m <= x"3d7d";
		r_c <= x"bc5f";
		wait for clk_period;
		x <= x"4964";
		y <= x"aa90";
		m <= x"7fd9";
		r_c <= x"d96a";
		wait for clk_period;
		x <= x"9f04";
		y <= x"454d";
		m <= x"e7f4";
		r_c <= x"ebb1";
		wait for clk_period;
		x <= x"5609";
		y <= x"d2a9";
		m <= x"3bfd";
		r_c <= x"e3bf";
		wait for clk_period;
		x <= x"fe37";
		y <= x"1a06";
		m <= x"270a";
		r_c <= x"f9fa";
		wait for clk_period;
		x <= x"5799";
		y <= x"c2f2";
		m <= x"246b";
		r_c <= x"18fa";
		wait for clk_period;
		x <= x"4b55";
		y <= x"03bc";
		m <= x"059b";
		r_c <= x"c4da";
		wait for clk_period;
		x <= x"1e47";
		y <= x"557e";
		m <= x"003d";
		r_c <= x"2d9a";
		wait for clk_period;
		x <= x"5e67";
		y <= x"f993";
		m <= x"f65d";
		r_c <= x"80c6";
		wait for clk_period;
		x <= x"5954";
		y <= x"6949";
		m <= x"9dee";
		r_c <= x"4ea3";
		wait for clk_period;
		x <= x"1e3f";
		y <= x"56c2";
		m <= x"0223";
		r_c <= x"c3f7";
		wait for clk_period;
		x <= x"ef19";
		y <= x"f4e7";
		m <= x"ef5b";
		r_c <= x"29de";
		wait for clk_period;
		x <= x"6944";
		y <= x"569d";
		m <= x"81ec";
		r_c <= x"2f96";
		wait for clk_period;
		x <= x"75cd";
		y <= x"5878";
		m <= x"84b4";
		r_c <= x"bb25";
		wait for clk_period;
		x <= x"b2b4";
		y <= x"f6ce";
		m <= x"7235";
		r_c <= x"3c63";
		wait for clk_period;
		x <= x"3fc9";
		y <= x"0a90";
		m <= x"8fd9";
		r_c <= x"92fe";
		wait for clk_period;
		x <= x"009e";
		y <= x"40c1";
		m <= x"e121";
		r_c <= x"e36c";
		wait for clk_period;
		x <= x"aa12";
		y <= x"1d37";
		m <= x"2bd2";
		r_c <= x"811f";
		wait for clk_period;
		x <= x"f132";
		y <= x"17b4";
		m <= x"238e";
		r_c <= x"a971";
		wait for clk_period;
		x <= x"6729";
		y <= x"c036";
		m <= x"a051";
		r_c <= x"1cb9";
		wait for clk_period;
		x <= x"3156";
		y <= x"b435";
		m <= x"0e50";
		r_c <= x"0e8d";
		wait for clk_period;
		x <= x"df5f";
		y <= x"ca76";
		m <= x"2fb2";
		r_c <= x"8b29";
		wait for clk_period;
		x <= x"c95a";
		y <= x"e78e";
		m <= x"db56";
		r_c <= x"4c6d";
		wait for clk_period;
		x <= x"28f5";
		y <= x"5071";
		m <= x"78aa";
		r_c <= x"308e";
		wait for clk_period;
		x <= x"2d32";
		y <= x"5104";
		m <= x"7986";
		r_c <= x"2fdb";
		wait for clk_period;
		x <= x"306f";
		y <= x"28ea";
		m <= x"bd5f";
		r_c <= x"4db5";
		wait for clk_period;
		x <= x"5e02";
		y <= x"ae05";
		m <= x"8507";
		r_c <= x"b28c";
		wait for clk_period;
		x <= x"3b7e";
		y <= x"bc2b";
		m <= x"9a41";
		r_c <= x"25b0";
		wait for clk_period;
		x <= x"f179";
		y <= x"3795";
		m <= x"5360";
		r_c <= x"61cd";
		wait for clk_period;
		x <= x"8fd1";
		y <= x"df3c";
		m <= x"ceda";
		r_c <= x"711a";
		wait for clk_period;
		x <= x"57f4";
		y <= x"2151";
		m <= x"b1fa";
		r_c <= x"396f";
		wait for clk_period;
		x <= x"9f22";
		y <= x"55f5";
		m <= x"00ef";
		r_c <= x"4b99";
		wait for clk_period;
		x <= x"e80b";
		y <= x"b18d";
		m <= x"0a54";
		r_c <= x"33f4";
		wait for clk_period;
		x <= x"98f4";
		y <= x"c5d4";
		m <= x"28bf";
		r_c <= x"bc9c";
		wait for clk_period;
		x <= x"ccb6";
		y <= x"2b06";
		m <= x"408a";
		r_c <= x"54fa";
		wait for clk_period;
		x <= x"adcf";
		y <= x"23f6";
		m <= x"b5f1";
		r_c <= x"83d0";
		wait for clk_period;
		x <= x"40f3";
		y <= x"2859";
		m <= x"3c85";
		r_c <= x"0c6b";
		wait for clk_period;
		x <= x"f98e";
		y <= x"df68";
		m <= x"4f1c";
		r_c <= x"561f";
		wait for clk_period;
		x <= x"636a";
		y <= x"b982";
		m <= x"1644";
		r_c <= x"b822";
		wait for clk_period;
		x <= x"004e";
		y <= x"3c9e";
		m <= x"daee";
		r_c <= x"867e";
		wait for clk_period;
		x <= x"f496";
		y <= x"1f6b";
		m <= x"af20";
		r_c <= x"5c39";
		wait for clk_period;
		x <= x"1268";
		y <= x"2c21";
		m <= x"c231";
		r_c <= x"c67f";
		wait for clk_period;
		x <= x"2e5a";
		y <= x"37b7";
		m <= x"5392";
		r_c <= x"8867";
		wait for clk_period;
		x <= x"c1d6";
		y <= x"e520";
		m <= x"57b0";
		r_c <= x"e4d1";
		wait for clk_period;
		x <= x"cd8f";
		y <= x"1d86";
		m <= x"ac4a";
		r_c <= x"a32b";
		wait for clk_period;
		x <= x"e4d2";
		y <= x"caef";
		m <= x"3066";
		r_c <= x"0f66";
		wait for clk_period;
		x <= x"36c6";
		y <= x"17dc";
		m <= x"23cb";
		r_c <= x"eeb6";
		wait for clk_period;
		x <= x"df4a";
		y <= x"d062";
		m <= x"3893";
		r_c <= x"936a";
		wait for clk_period;
		x <= x"eace";
		y <= x"e7c4";
		m <= x"5ba7";
		r_c <= x"cbe2";
		wait for clk_period;
		x <= x"1819";
		y <= x"f6be";
		m <= x"f21e";
		r_c <= x"580f";
		wait for clk_period;
		x <= x"02ad";
		y <= x"0b73";
		m <= x"912d";
		r_c <= x"588e";
		wait for clk_period;
		x <= x"b244";
		y <= x"5a01";
		m <= x"0701";
		r_c <= x"6b43";
		wait for clk_period;
		x <= x"fafd";
		y <= x"942b";
		m <= x"5e41";
		r_c <= x"c35e";
		wait for clk_period;
		x <= x"4145";
		y <= x"ba77";
		m <= x"17b3";
		r_c <= x"c5d1";
		wait for clk_period;
		x <= x"cf69";
		y <= x"745c";
		m <= x"2e8b";
		r_c <= x"a3a1";
		wait for clk_period;
		x <= x"8061";
		y <= x"ee91";
		m <= x"e5da";
		r_c <= x"b3d4";
		wait for clk_period;
		x <= x"3c6c";
		y <= x"ebd9";
		m <= x"e1c6";
		r_c <= x"5780";
		wait for clk_period;
		x <= x"c52e";
		y <= x"9553";
		m <= x"dffd";
		r_c <= x"8e09";
		wait for clk_period;
		x <= x"4bb5";
		y <= x"ff64";
		m <= x"7f16";
		r_c <= x"051d";
		wait for clk_period;
		x <= x"c6f4";
		y <= x"98a2";
		m <= x"e4f4";
		r_c <= x"0987";
		wait for clk_period;
		x <= x"a2f9";
		y <= x"1382";
		m <= x"1d43";
		r_c <= x"4fc6";
		wait for clk_period;
		x <= x"48e9";
		y <= x"e7e4";
		m <= x"dbd6";
		r_c <= x"2c45";
		wait for clk_period;
		x <= x"6b21";
		y <= x"503b";
		m <= x"7859";
		r_c <= x"4d3c";
		wait for clk_period;
		x <= x"38b1";
		y <= x"c898";
		m <= x"ace4";
		r_c <= x"8473";
		wait for clk_period;
		x <= x"9640";
		y <= x"aa95";
		m <= x"7fe0";
		r_c <= x"ac49";
		wait for clk_period;
		x <= x"f044";
		y <= x"ead5";
		m <= x"e040";
		r_c <= x"9d68";
		wait for clk_period;
		x <= x"6099";
		y <= x"3dcd";
		m <= x"dcb4";
		r_c <= x"2e2f";
		wait for clk_period;
		x <= x"e375";
		y <= x"8edf";
		m <= x"564e";
		r_c <= x"58ee";
		wait for clk_period;
		x <= x"799f";
		y <= x"e88d";
		m <= x"dcd4";
		r_c <= x"b2b7";
		wait for clk_period;
		x <= x"b555";
		y <= x"ecdf";
		m <= x"e34f";
		r_c <= x"80f9";
		wait for clk_period;
		x <= x"e474";
		y <= x"a343";
		m <= x"74e5";
		r_c <= x"c8fa";
		wait for clk_period;
		x <= x"e671";
		y <= x"23f7";
		m <= x"35f3";
		r_c <= x"a7a8";
		wait for clk_period;
		x <= x"9545";
		y <= x"2314";
		m <= x"349e";
		r_c <= x"5dad";
		wait for clk_period;
		x <= x"e3f5";
		y <= x"a034";
		m <= x"704e";
		r_c <= x"b4f0";
		wait for clk_period;
		x <= x"f191";
		y <= x"16a5";
		m <= x"a1f8";
		r_c <= x"9466";
		wait for clk_period;
		x <= x"944e";
		y <= x"9883";
		m <= x"e4c4";
		r_c <= x"e3f8";
		wait for clk_period;
		x <= x"5cd6";
		y <= x"366c";
		m <= x"d1a2";
		r_c <= x"c095";
		wait for clk_period;
		x <= x"2b47";
		y <= x"052d";
		m <= x"07c3";
		r_c <= x"d244";
		wait for clk_period;
		x <= x"fc9b";
		y <= x"2026";
		m <= x"3039";
		r_c <= x"c724";
		wait for clk_period;
		x <= x"09e3";
		y <= x"1f1e";
		m <= x"aead";
		r_c <= x"2163";
		wait for clk_period;
		x <= x"a120";
		y <= x"3351";
		m <= x"4cf9";
		r_c <= x"19d8";
		wait for clk_period;
		x <= x"132a";
		y <= x"2dc6";
		m <= x"c4a9";
		r_c <= x"42b9";
		wait for clk_period;
		x <= x"729f";
		y <= x"c915";
		m <= x"ad9f";
		r_c <= x"7468";
		wait for clk_period;
		x <= x"1566";
		y <= x"88fd";
		m <= x"cd7c";
		r_c <= x"d353";
		wait for clk_period;
		x <= x"f5f3";
		y <= x"bab2";
		m <= x"180b";
		r_c <= x"55b8";
		wait for clk_period;
		x <= x"95ad";
		y <= x"5306";
		m <= x"7c8a";
		r_c <= x"a27f";
		wait for clk_period;
		x <= x"8f5c";
		y <= x"0768";
		m <= x"8b1c";
		r_c <= x"203c";
		wait for clk_period;
		x <= x"d322";
		y <= x"1b23";
		m <= x"28b4";
		r_c <= x"ab11";
		wait for clk_period;
		x <= x"06f2";
		y <= x"4eac";
		m <= x"f602";
		r_c <= x"0a4a";
		wait for clk_period;
		x <= x"e023";
		y <= x"6b6f";
		m <= x"a126";
		r_c <= x"542e";
		wait for clk_period;
		x <= x"b7e5";
		y <= x"44aa";
		m <= x"e6ff";
		r_c <= x"8677";
		wait for clk_period;
		x <= x"1793";
		y <= x"a611";
		m <= x"7919";
		r_c <= x"acb2";
		wait for clk_period;
		x <= x"fd1f";
		y <= x"04a5";
		m <= x"86f8";
		r_c <= x"b221";
		wait for clk_period;
		x <= x"7f48";
		y <= x"65b1";
		m <= x"1889";
		r_c <= x"5497";
		wait for clk_period;
		x <= x"0225";
		y <= x"537f";
		m <= x"7d3f";
		r_c <= x"707a";
		wait for clk_period;
		x <= x"00f0";
		y <= x"9b4a";
		m <= x"e8ef";
		r_c <= x"8324";	
		wait for clk_period;
		valid_in <= '0';

--valid_in <='0';


      wait;
   end process;

END;
